package ve_package;

`include "ve_base_unit.svh"
`include "ve_operands.svh"
`include "ve_result.svh"
`include "ve_rst_bfm.svh"
`include "ve_data_in_generator.svh"
`include "ve_data_in_bfm.svh"
`include "ve_data_out_generator.svh"
`include "ve_data_out_bfm.svh"
`include "ve_environment.svh"

endpackage
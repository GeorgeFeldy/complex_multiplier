library verilog;
use verilog.vl_types.all;
entity complex_multiplier_test is
end complex_multiplier_test;
